--------------------------------------------------------------------------------
-- Project : PROJECTNAME
-- Author : Donald MacIntyre - djm4912
-- Date : 4/8/2018
-- File : lms.vhd
--------------------------------------------------------------------------------
-- Description :
--------------------------------------------------------------------------------
-- $Log$
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

use work.lms_pkg.all;

entity lms is
    Port (
        clk         : in std_logic;
        rst         : in std_logic;
        in_valid    : in std_logic;
        xin         : in signed(15 downto 0);
        expected    : in signed(15 downto 0);
        out_valid   : out std_logic
    );
end lms;

architecture behav of lms is

--------------------------------------------------------------------------------
-- Signal Declarations
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Component Declarations
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------

begin

end behav;