library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work ;

package lms_pkg is

end package lms_pkg;
